module or_gate_8(c,i1,i2,i3,i4,i5,i6,i7,i8);
output c;
input i1,i2,i3,i4,i5,i6,i7,i8;
wire w1,w2,w3,w4,w5,w6,w7,w8,w9,w10;
wire w11,w12,w13,w14,w15,w16,w17,w18,w19,w20;
nand(w1,i1,i1);
nand(w2,i2,i2);
nand(w3,w1,w2);
nand(w4,i3,i3);
nand(w5,i4,i4);
nand(w6,w4,w5);
nand(w7,i5,i5);
nand(w8,i6,i6);
nand(w9,w7,w8);
nand(w10,i7,i7);
nand(w11,i8,i8);
nand(w12,w10,w11);
nand(w13,w3,w3);
nand(w14,w6,w6);
nand(w15,w13,w14);
nand(w16,w9,w9);
nand(w17,w12,w12);
nand(w18,w16,w17);
nand(w19,w15,w15);
nand(w20,w18,w18);
nand(c,w19,w20);
endmodule
