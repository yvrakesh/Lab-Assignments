
module not_gate(b,a);
output b;
input a;
nand(b,a,a);
endmodule