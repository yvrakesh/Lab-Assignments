module mux_1_2(y,s,a,b);
output y;
input s,a,b;
wire p,q,r;
nand(p,s,s);
nand(q,p,a);
nand(r,s,b);
nand(y,q,r);
endmodule
